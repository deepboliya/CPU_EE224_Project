
library ieee;
use ieee.std_logic_1164.all;

entity MUX_1_TO_5 is
    port(
        i: in std_logic_vector(15 downto 0);
        D0,D1,D2,D3,D4: out std_logic_vector(15 downto 0);
        S: in std_logic_vector(2 downto 0)
         );
end MUX_1_TO_5;
architecture Struct of MUX_1_to_5 is

begin
	process( i,S )
	begin
	 case s is
		when"000" =>
		d0<=i;
		d1<="0000000000000000";
		d2<="0000000000000000";
		d3<="0000000000000000";
		d4<="0000000000000000";
		when "001"=>
		d1<=i;
		d0<="0000000000000000";
		d2<="0000000000000000";
		d3<="0000000000000000";
		d4<="0000000000000000";
		when "010" =>
		d2<=i;
		d1<="0000000000000000";
		d3<="0000000000000000";
		d4<="0000000000000000";
		d0<="0000000000000000";
		when "011" =>
		d3<=i;
		d1<="0000000000000000";
		d0<="0000000000000000";
		d2<="0000000000000000";
		d4<="0000000000000000";
		when "100" =>
		d4<=i;
		d0<="0000000000000000";
		d1<="0000000000000000";
		d3<="0000000000000000";
		d2<="0000000000000000";
		
		when others=>
		d2<="0000000000000000";
		d0<="0000000000000000";
		d1<="0000000000000000";
		d3<="0000000000000000";
		d4<="0000000000000000";
		end case;
	end process; 
	
end Struct;